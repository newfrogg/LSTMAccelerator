package accel_pkg;
    
    // Accelerator constants
    parameter int unsigned ELEMENT_BITS = 32;

    
endpackage