`timescale 1ps / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/07/2024 03:22:42 PM
// Design Name: 
// Module Name: tb_tanh
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_tanh();
    
    reg     [31:0] data_in;
    wire    [7:0] data_out;
    tanh t0 ( .data_in(data_in), .data_out(data_out) );
    int k = 0;
    initial begin
        data_in = 32'h80000006;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h90041d37;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h9973a50f;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'ha56ceffc;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'ha9bab234;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'had623a06;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hb0900e11;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hb360eb90;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hb5e87484;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hb834ab38;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hba4fe888;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hbc420896;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hbe1127d5;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hbfc21ebc;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hc158d57d;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hc2d87e59;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hc443bf3e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hc59cd028;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hc6e591ae;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hc81f9e17;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hc94c566f;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hca6cecb4;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hcb826bd9;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hcc8dbe2b;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hcd8fb26a;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hce88fff8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hcf7a4a3a;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hd064236c;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hd1470ef1;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hd2238346;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hd2f9eba8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hd3caa973;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hd4961554;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hd55c8048;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hd61e347b;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hd6db7607;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hd7948399;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hd8499706;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hd8fae5c2;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hd9a8a153;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hda52f7b1;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hdafa139d;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hdb9e1cea;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hdc3f38c3;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hdcdd89e8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hdd7930de;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hde124c25;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hdea8f861;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hdf3d507e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hdfcf6dd7;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he05f6852;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he0ed567f;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he1794daf;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he203620f;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he28ba6ba;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he3122dce;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he397087e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he41a4721;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he49bf942;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he51c2dad;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he59af27c;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he6185523;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he6946278;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he70f26c2;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he788adbb;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he80102a0;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he8783032;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he8ee40c1;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he9633e33;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he9d73209;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hea4a2562;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'heabc2109;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'heb2d2d6e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'heb9d52b5;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hec0c98b6;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hec7b0701;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hece8a4e1;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hed557964;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hedc18b59;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hee2ce157;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hee9781bd;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hef0172b7;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hef6aba42;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hefd35e29;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf03b640d;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf0a2d166;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf109ab82;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf16ff78a;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf1d5ba83;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf23af952;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf29fb8b7;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf303fd58;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf367cbba;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf3cb2849;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf42e1755;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf4909d15;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf4f2bda7;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf5547d16;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf5b5df53;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf616e83e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf6779ba2;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf6d7fd37;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf73810a6;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf797d986;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf7f75b5d;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf85699a6;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf8b597ca;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf9145929;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf972e114;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf9d132d0;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hfa2f519b;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hfa8d40a4;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hfaeb0314;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hfb489c0a;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hfba60e9e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hfc035ddf;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hfc608cd6;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hfcbd9e86;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hfd1a95ec;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hfd777601;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hfdd441b8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hfe30fc01;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hfe8da7c9;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hfeea47fa;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hff46df7b;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hffa37133;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h6;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h5c8ed7;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hb9208f;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h115b810;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h1725841;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h1cf0409;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h22bbe52;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h2888a09;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h2e56a1e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h3426184;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h39f7334;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h3fca22b;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h459f16c;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h4b76400;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h514fcf6;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h572bf66;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h5d0ae6f;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h62ecd3a;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h68d1ef6;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h6eba6e1;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h74a6840;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h7a96664;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h808a4ad;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h8682684;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h8c7ef64;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h92802d3;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h9886468;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h9e917cc;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'ha4a20b7;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'haab82f4;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hb0d4263;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hb6f62f5;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hbd1e8b5;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hc34d7c1;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hc983450;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hcfc02b2;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hd604753;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hdc506b8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he2a4587;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'he900880;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hef65488;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hf5d2ea4;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'hfc49bfd;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h102ca1e1;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h109545c8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h10fe8d53;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h11687e4d;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h11d31eb3;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h123e74b1;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h12aa86a6;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h13175b29;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h1384f909;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h13f36754;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h1462ad55;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h14d2d29c;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h1543df01;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h15b5daa8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h1628ce01;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h169cc1d7;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h1711bf49;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h1787cfd8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h17fefd6a;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h1877524f;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h18f0d948;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h196b9d92;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h19e7aae7;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h1a650d8e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h1ae3d25d;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h1b6406c8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h1be5b8e9;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h1c68f78c;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h1cedd23c;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h1d745950;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h1dfc9dfb;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h1e86b25b;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h1f12a98b;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h1fa097b8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h20309233;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h20c2af8c;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h215707a9;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h21edb3e5;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h2286cf2c;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h23227622;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h23c0c747;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h2461e320;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h2505ec6d;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h25ad0859;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h26575eb7;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h27051a48;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h27b66904;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h286b7c71;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h29248a03;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h29e1cb8f;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h2aa37fc2;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h2b69eab6;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h2c355697;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h2d061462;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h2ddc7cc4;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h2eb8f119;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h2f9bdc9e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h3085b5d0;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h31770012;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h32704da0;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h337241df;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h347d9431;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h35931356;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h36b3a99b;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h37e061f3;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h391a6e5c;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h3a632fe2;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h3bbc40cc;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h3d2781b1;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h3ea72a8d;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h403de14e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h41eed835;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h43bdf774;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h45b01782;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h47cb54d2;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h4a178b86;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h4c9f147a;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h4f6ff1f9;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h529dc604;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h56454dd6;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h5a93100e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h5fd19313;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h668c5afb;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
        data_in = 32'h6ffbe2d3;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k = k+1;
    end
    
endmodule

