`timescale 1ps / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/08/2024 08:38:40 AM
// Design Name: 
// Module Name: tb_sigmoid
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_sigmoid();
    reg     [31:0] data_in;
    wire    [7:0] data_out;
    sigmoid s0 ( .data_in(data_in), .data_out(data_out) );
    int k = 0;
    initial begin
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h81922537;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h9163fffe;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h9ab5ebf3;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'ha15b95ef;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'ha689a465;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'haac9e593;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hae65f605;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hb189d09d;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hb451d866;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hb6d171c5;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hb916730d;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hbb2b14a3;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hbd1719fe;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hbee08c64;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hc08c3516;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hc21df005;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hc398e569;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hc4ffb2e1;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hc6548972;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hc79943d0;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hc8cf773a;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hc9f88067;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hcb158d95;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hcc27a673;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hcd2fb26d;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hce2e7dbb;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hcf24bd7f;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hd013131f;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hd0fa0f09;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hd1da3306;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hd2b3f41f;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hd387bc40;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hd455eb94;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hd51ed9b0;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hd5e2d695;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hd6a22b85;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hd75d1bc5;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hd813e53e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hd8c6c10d;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hd975e401;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hda217f03;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hdac9bf7b;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hdb6ecfa4;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hdc10d6d5;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hdcaff9c3;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hdd4c5ac1;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hdde619ef;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hde7d556e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hdf122985;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hdfa4b0ce;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he0350454;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he0c33bb3;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he14f6d32;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he1d9ade1;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he26211ac;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he2e8ab74;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he36d8d1d;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he3f0c7a3;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he4726b2c;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he4f28712;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he57129f1;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he5ee61b9;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he66a3bb1;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he6e4c48a;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he75e0861;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he7d612ce;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he84ceee9;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he8c2a752;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he937463a;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he9aad566;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hea1d5e39;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hea8ee9b8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'heaff808f;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'heb6f2b17;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hebddf158;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hec4bdb13;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hecb8efbe;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hed253690;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hed90b680;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hedfb7646;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hee657c66;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'heececf2b;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hef3774ae;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hef9f72d8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf006cf62;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf06d8fdd;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf0d3b9ae;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf1395214;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf19e5e27;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf202e2dc;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf266e509;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf2ca6960;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf32d7477;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf3900ac6;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf3f230ab;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf453ea68;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf4b53c26;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf51629fa;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf576b7de;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf5d6e9b9;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf636c35e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf696488c;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf6f57cf1;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf7546429;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf7b301c0;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf8115932;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf86f6dee;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf8cd4353;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf92adcb7;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf9883d5f;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf9e56889;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hfa426164;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hfa9f2b1a;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hfafbc8c8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hfb583d84;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hfbb48c5b;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hfc10b854;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hfc6cc46e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hfcc8b3a2;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hfd2488e6;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hfd804727;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hfddbf150;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hfe378a49;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hfe9314f4;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hfeee9433;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hff4a0ae5;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hffa57be6;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hea14;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h5c5848;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hb7c95f;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h1134036;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h16ebfa8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h1ca4a96;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h225e3df;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h2818e68;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h2dd4d18;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h33922d8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h395129a;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h3f11f4f;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h44d4bf3;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h4a99b84;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h506110a;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h562af92;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h5bf7a31;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h61c7406;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h679a03a;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h6d701fc;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h7349c8b;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h792732c;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h7f08935;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h84ee206;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h8ad810d;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h90c69c7;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h96b9fc1;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h9cb2696;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'ha2b01f5;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'ha8b359e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'haebc563;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hb4cb52c;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hbae08f5;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hc0fc4d1;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hc71ecea;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hcd48584;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hd3792fd;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hd9b19cd;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hdff1e8a;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'he63a5e8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hec8b4bd;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf2e4ffe;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hf947cc5;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'hffb4051;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h1062a00a;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h10caa17d;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h11334a69;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h119ca0b4;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h1206aa7b;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h12716e09;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h12dcf1e1;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h13493cc0;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h13b6559c;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h142443ac;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h14930e6b;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h1502bd98;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h1573593e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h15e4e9b8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h165777b4;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h16cb0c37;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h173fb0a7;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h17b56ecc;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h182c50d8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h18a4616e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h191daba7;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h19983b1f;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h1a141bf6;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h1a915adf;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h1b100525;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h1b9028ba;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h1c11d440;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h1c951714;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h1d1a015f;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h1da0a422;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h1e291147;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h1eb35bb3;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h1f3f9757;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h1fcdd94a;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h205e37da;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h20f0caaa;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h2185aacc;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h221cf2e2;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h22b6bf3d;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h23532e07;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h23f25f6b;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h249475c8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h253995df;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h25e1e717;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h268d93b8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h273cc93c;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h27efb8a1;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h28a696c8;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h29619ce7;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h2a210900;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h2ae51e75;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h2bae26ab;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h2c7c71c4;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h2d505780;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h2e2a3839;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h2f0a7e10;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h2ff19e4c;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h30e01af9;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h31d684d9;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h32d57dae;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h33ddbb08;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h34f0099e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h360d5175;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h37369aef;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h386d1524;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h39b21dcf;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h3b074b72;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h3c6e7a4c;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h3de9dd4f;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h3f7c148e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h41284b66;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h42f261e6;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h44df26cc;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h46f4aad9;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h493abbfd;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h4bbba1bf;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h4e854925;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h51ab3a3e;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h554a1386;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h598e3ae0;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h5ec222d6;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h65718cfb;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h6ed6f9c7;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
        data_in = 32'h7ee358a0;
        #10;
        $display("tests = %d, time = %0t, data_in = %h (hex), data_out = %b ", k, $time, data_in, data_out);
        k=k+1;
    end
endmodule

