module accel_top import accel_pkg::*; #(

) (
    input logic clk_i,
    input logic rst_ni,
    input logic en_weight_i,
    input logic en_bias_i,

    output logic predicted_valid_o
);

endmodule 